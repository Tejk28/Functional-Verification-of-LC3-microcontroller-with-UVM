package decode_env_pkg;

import uvm_pkg::*;
import uvmf_base_pkg::*;
import decode_in_pkg::*;
import decode_in_pkg_hdl::*;
import decode_out_pkg::*;
import decode_out_pkg_hdl::*;
`include "uvm_macros.svh"
`include "src/lc3_prediction_typedefs.svh"
`include "src/decode_model.svh"
`include "src/decode_env_configuration.svh"
`include "src/decode_scoreboard.svh"
`include "src/decode_predictor.svh"
`include "src/decode_environment.svh"

endpackage
