package lc3_prediction_pkg;

   import uvm_pkg::*;
   `include "src/lc3_prediction_typedefs.svh"
   `include "src/decode_model.svh"

endpackage
